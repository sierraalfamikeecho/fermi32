module memory #(
    parameter WORDS = 128,
    parameter mem_init = ""
)
(
    input logic clk,
    input logic [31:0] address,
    input logic [31:0] write_data,
    input logic [3:0] byte_enable,
    input logic write_enable,
    input logic nrst,

    output logic [31:0] read_data
);

reg [31:0] mem [0:WORDS-1];

initial begin
    if (mem_init != "") begin
        $readmemh(mem_init, mem);
    end
end

always @(posedge clk) begin
    if (nrst == 1'b0) begin
        for (int i  = 0; i < WORDS; i++) begin
            mem[i] <= 32'b0;
        end
        for (int i = 0; i < WORDS; i++) begin
            mem[i] <= 32'b0;
        end
    end else begin
        if(write_enable) begin
            if(address[1:0] != 2'b00) begin
                $display("misaligned write  at address %h", address);
            end else begin
                for (int i = 0; i < 4; i++) begin
                    if (byte_enable[i]) begin
                        mem[address[31:2]][(i*8)+:8] <= write_data[(i*8)+:8];
                    end
                end
            end
        end
    end
end

always_comb begin
    read_data = mem[address[31:2]];
end

endmodule
